// Convert a nine segment signal to a 3x3 anode common LED pins (6 pins)
module nine_segment_to_six_pin(
	input bit [8:0] segments,
	output logic [5:0] pins);
endmodule